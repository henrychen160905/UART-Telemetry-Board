module transmitter(
    input logic clk,
    input logic rst,
    input logic data_in,
    input logic start_signal,
    output logic transmit_wire,
    output logic state_busy
)
endmodule
