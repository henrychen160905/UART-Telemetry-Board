module transmitter(input logic clk, output logic tx);
    assign tx = clk;
endmodule
