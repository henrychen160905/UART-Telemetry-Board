module receiver(input logic rx, output logic valid);
    assign valid = rx;
endmodule

